module FoodLogic(
	input clk,
	input rst,
	output reg [7:0] x,
	output reg [6:0] y,
	output plotEn

);

endmodule