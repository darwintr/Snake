module drawBlack(
		input clk
	)