
module highscoreSystem(
	input clk,
	input rst,
	input increment,
	output reg [3:0] hex2_out, hex3_out
);
	reg [12:0] curr_score;
	

endmodule